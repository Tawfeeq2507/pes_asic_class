vim opt_check.v
``` verilog
module opt_check (input a , input b , output y);
        assign y = a?b:0;
endmodule
```
